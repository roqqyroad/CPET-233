--Name: Rachel DuBois
--Section: 02
--Lab: 02
--Assignment: Lab Eight - Counter
--Summary: Keeps count of how many times delay unit has been activated. 

--libraries
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

--START OF ENTITY

--END OF ENTITY

--START OF ARCHITECTURE

--END OF ARCHITECTURE