--Name: Rachel DuBois
--Section: 02
--Lab: 02
--Assignment: Homework Six - Question Five

--libraries
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;