--Name: Rachel DuBois
--Section: 02
--Lab: 02
--Assignment: Lab Six - Is Negative

entity is_neg is
    port(

    );
end is_neg;

architecture model of is_neg is

    begin
    
end model;