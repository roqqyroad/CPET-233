--Name: Rachel DuBois
--Section: 02
--Lab: 02
--Assignment: Homework Five - Question Two

entity question_two is
    port(

    );
end question_two;

architecture model of question_two is

begin

end model;

