--Name: Rachel DuBois
--Section: 02
--Lab: 02
--Assignment: Lab Six - Absolute Value

entity abs is
    port(

    );
end abs;

architecture model of abs is

begin

end model;

