--Name: Rachel DuBois
--Section: 02
--Lab: 02
--Assignment: Lab Six - Convert To Constant

entity convert_to_constant is
    port(

    );
end convert_to_constant;

architecture model of convert_to_constant is

    begin
        
end model;